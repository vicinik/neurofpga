library ieee;
use ieee.std_logic_1164;
use ieee.math_real;
use work.Global.all;

entity Layer is

end entity;

architecture Bhv of Layer is
	
begin
	
end architecture;