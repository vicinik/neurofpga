library ieee;
use ieee.std_logic_1164;
use ieee.math_real;
use work.Global.all;

entity Neuron is

end entity;

architecture Bhv of Neuron is
	
begin
	
end architecture;