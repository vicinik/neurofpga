library ieee;
use ieee.std_logic_1164;
use ieee.math_real;
use work.Global.all;

entity Net is

end entity;

architecture Bhv of Net is
	
begin
	
end architecture;